magic
tech sky130A
timestamp 1731942359
<< error_p >>
rect 95 -375 97 -350
<< nwell >>
rect -100 -350 200 65
<< nmos >>
rect 40 -500 55 -400
<< pmos >>
rect 40 -305 55 -95
<< ndiff >>
rect -5 -410 40 -400
rect -5 -490 5 -410
rect 25 -490 40 -410
rect -5 -500 40 -490
rect 55 -410 100 -400
rect 55 -490 70 -410
rect 90 -490 100 -410
rect 55 -500 100 -490
<< pdiff >>
rect -10 -105 40 -95
rect -10 -295 0 -105
rect 25 -295 40 -105
rect -10 -305 40 -295
rect 55 -105 105 -95
rect 55 -295 70 -105
rect 95 -295 105 -105
rect 55 -305 105 -295
<< ndiffc >>
rect 5 -490 25 -410
rect 70 -490 90 -410
<< pdiffc >>
rect 0 -295 25 -105
rect 70 -295 95 -105
<< psubdiff >>
rect -10 -550 105 -535
rect -10 -570 5 -550
rect 90 -570 105 -550
rect -10 -585 105 -570
<< nsubdiff >>
rect -30 15 125 30
rect -30 -15 -15 15
rect 110 -15 125 15
rect -30 -30 125 -15
<< psubdiffcont >>
rect 5 -570 90 -550
<< nsubdiffcont >>
rect -15 -15 110 15
<< poly >>
rect 40 -95 55 -50
rect 40 -335 55 -305
rect -10 -380 55 -335
rect 40 -400 55 -380
rect 40 -525 55 -500
<< locali >>
rect -30 20 125 30
rect -30 15 20 20
rect 65 15 125 20
rect -30 -15 -15 15
rect 110 -15 125 15
rect -30 -20 20 -15
rect 65 -20 125 -15
rect -30 -30 125 -20
rect -10 -105 35 -30
rect -10 -295 0 -105
rect 25 -295 35 -105
rect -10 -305 35 -295
rect 60 -105 105 -95
rect 60 -295 70 -105
rect 95 -295 105 -105
rect 60 -305 105 -295
rect 60 -330 100 -305
rect -10 -345 30 -335
rect -10 -370 0 -345
rect 20 -370 30 -345
rect -10 -380 30 -370
rect 60 -350 120 -330
rect 60 -375 80 -350
rect 95 -375 120 -350
rect 60 -390 120 -375
rect -5 -410 35 -400
rect -5 -490 5 -410
rect 25 -475 35 -410
rect 60 -410 100 -390
rect 25 -490 40 -475
rect -5 -540 40 -490
rect 60 -490 70 -410
rect 90 -490 100 -410
rect 60 -500 100 -490
rect -5 -545 100 -540
rect -5 -550 25 -545
rect 55 -550 100 -545
rect -5 -570 5 -550
rect 90 -570 100 -550
rect -5 -575 25 -570
rect 55 -575 100 -570
rect -5 -580 100 -575
rect -5 -585 40 -580
<< viali >>
rect 20 15 65 20
rect 20 -15 65 15
rect 20 -20 65 -15
rect 0 -370 20 -345
rect 80 -375 95 -350
rect 25 -550 55 -545
rect 25 -570 55 -550
rect 25 -575 55 -570
<< metal1 >>
rect -295 20 430 30
rect -295 -20 20 20
rect 65 -20 430 20
rect -295 -30 430 -20
rect -200 -345 30 -335
rect -200 -370 0 -345
rect 20 -370 30 -345
rect -200 -380 30 -370
rect 60 -350 425 -330
rect 60 -375 80 -350
rect 95 -375 425 -350
rect 60 -390 425 -375
rect -280 -545 430 -535
rect -280 -575 25 -545
rect 55 -575 430 -545
rect -280 -590 430 -575
<< end >>
